// Nios.v

// Generated using ACDS version 13.1 162 at 2018.10.22.15:29:04

`timescale 1 ps / 1 ps
module Nios (
		input  wire        clk_clk,                                     //                              clk.clk
		input  wire        pushbutton2_external_connection_export,      //  pushbutton2_external_connection.export
		output wire        led_1_external_connection_export,            //        led_1_external_connection.export
		output wire        led_2_external_connection_export,            //        led_2_external_connection.export
		output wire        led_3_external_connection_export,            //        led_3_external_connection.export
		output wire        led_4_external_connection_export,            //        led_4_external_connection.export
		output wire        led_5_external_connection_export,            //        led_5_external_connection.export
		input  wire        pushbutton_1_external_connection_export,     // pushbutton_1_external_connection.export
		input  wire        dip_0_external_connection_export,            //        dip_0_external_connection.export
		input  wire        dip_1_external_connection_export,            //        dip_1_external_connection.export
		input  wire        dip_2_external_connection_export,            //        dip_2_external_connection.export
		input  wire        dip_3_external_connection_export,            //        dip_3_external_connection.export
		output wire        lcd_0_conduit_end_rs,                        //                lcd_0_conduit_end.rs
		output wire        lcd_0_conduit_end_rw,                        //                                 .rw
		output wire        lcd_0_conduit_end_en,                        //                                 .en
		output wire [7:0]  lcd_0_conduit_end_db,                        //                                 .db
		input  wire        eth_tse_0_mac_status_connection_set_10,      //  eth_tse_0_mac_status_connection.set_10
		input  wire        eth_tse_0_mac_status_connection_set_1000,    //                                 .set_1000
		output wire        eth_tse_0_mac_status_connection_eth_mode,    //                                 .eth_mode
		output wire        eth_tse_0_mac_status_connection_ena_10,      //                                 .ena_10
		input  wire [7:0]  eth_tse_0_mac_gmii_connection_gmii_rx_d,     //    eth_tse_0_mac_gmii_connection.gmii_rx_d
		input  wire        eth_tse_0_mac_gmii_connection_gmii_rx_dv,    //                                 .gmii_rx_dv
		input  wire        eth_tse_0_mac_gmii_connection_gmii_rx_err,   //                                 .gmii_rx_err
		output wire [7:0]  eth_tse_0_mac_gmii_connection_gmii_tx_d,     //                                 .gmii_tx_d
		output wire        eth_tse_0_mac_gmii_connection_gmii_tx_en,    //                                 .gmii_tx_en
		output wire        eth_tse_0_mac_gmii_connection_gmii_tx_err,   //                                 .gmii_tx_err
		input  wire [3:0]  eth_tse_0_mac_mii_connection_mii_rx_d,       //     eth_tse_0_mac_mii_connection.mii_rx_d
		input  wire        eth_tse_0_mac_mii_connection_mii_rx_dv,      //                                 .mii_rx_dv
		input  wire        eth_tse_0_mac_mii_connection_mii_rx_err,     //                                 .mii_rx_err
		output wire [3:0]  eth_tse_0_mac_mii_connection_mii_tx_d,       //                                 .mii_tx_d
		output wire        eth_tse_0_mac_mii_connection_mii_tx_en,      //                                 .mii_tx_en
		output wire        eth_tse_0_mac_mii_connection_mii_tx_err,     //                                 .mii_tx_err
		input  wire        eth_tse_0_mac_mii_connection_mii_crs,        //                                 .mii_crs
		input  wire        eth_tse_0_mac_mii_connection_mii_col,        //                                 .mii_col
		output wire        eth_tse_0_mac_misc_connection_magic_wakeup,  //    eth_tse_0_mac_misc_connection.magic_wakeup
		input  wire        eth_tse_0_mac_misc_connection_magic_sleep_n, //                                 .magic_sleep_n
		input  wire        eth_tse_0_mac_misc_connection_ff_tx_crc_fwd, //                                 .ff_tx_crc_fwd
		output wire        eth_tse_0_mac_misc_connection_ff_tx_septy,   //                                 .ff_tx_septy
		output wire        eth_tse_0_mac_misc_connection_tx_ff_uflow,   //                                 .tx_ff_uflow
		output wire        eth_tse_0_mac_misc_connection_ff_tx_a_full,  //                                 .ff_tx_a_full
		output wire        eth_tse_0_mac_misc_connection_ff_tx_a_empty, //                                 .ff_tx_a_empty
		output wire [17:0] eth_tse_0_mac_misc_connection_rx_err_stat,   //                                 .rx_err_stat
		output wire [3:0]  eth_tse_0_mac_misc_connection_rx_frm_type,   //                                 .rx_frm_type
		output wire        eth_tse_0_mac_misc_connection_ff_rx_dsav,    //                                 .ff_rx_dsav
		output wire        eth_tse_0_mac_misc_connection_ff_rx_a_full,  //                                 .ff_rx_a_full
		output wire        eth_tse_0_mac_misc_connection_ff_rx_a_empty  //                                 .ff_rx_a_empty
	);

	wire         nios_jtag_debug_module_reset_reset;                                      // Nios:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire  [31:0] nios_custom_instruction_master_result;                                   // Nios_custom_instruction_master_translator:ci_slave_result -> Nios:E_ci_result
	wire   [4:0] nios_custom_instruction_master_b;                                        // Nios:D_ci_b -> Nios_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_c;                                        // Nios:D_ci_c -> Nios_custom_instruction_master_translator:ci_slave_c
	wire         nios_custom_instruction_master_done;                                     // Nios_custom_instruction_master_translator:ci_slave_multi_done -> Nios:E_ci_multi_done
	wire         nios_custom_instruction_master_clk_en;                                   // Nios:E_ci_multi_clk_en -> Nios_custom_instruction_master_translator:ci_slave_multi_clken
	wire   [4:0] nios_custom_instruction_master_a;                                        // Nios:D_ci_a -> Nios_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] nios_custom_instruction_master_n;                                        // Nios:D_ci_n -> Nios_custom_instruction_master_translator:ci_slave_n
	wire         nios_custom_instruction_master_writerc;                                  // Nios:D_ci_writerc -> Nios_custom_instruction_master_translator:ci_slave_writerc
	wire         nios_custom_instruction_master_clk;                                      // Nios:E_ci_multi_clock -> Nios_custom_instruction_master_translator:ci_slave_multi_clk
	wire         nios_custom_instruction_master_reset_req;                                // Nios:E_ci_multi_reset_req -> Nios_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios_custom_instruction_master_start;                                    // Nios:E_ci_multi_start -> Nios_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] nios_custom_instruction_master_dataa;                                    // Nios:E_ci_dataa -> Nios_custom_instruction_master_translator:ci_slave_dataa
	wire         nios_custom_instruction_master_readra;                                   // Nios:D_ci_readra -> Nios_custom_instruction_master_translator:ci_slave_readra
	wire         nios_custom_instruction_master_reset;                                    // Nios:E_ci_multi_reset -> Nios_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] nios_custom_instruction_master_datab;                                    // Nios:E_ci_datab -> Nios_custom_instruction_master_translator:ci_slave_datab
	wire         nios_custom_instruction_master_readrb;                                   // Nios:D_ci_readrb -> Nios_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_result;        // Nios_custom_instruction_master_multi_xconnect:ci_slave_result -> Nios_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_b;             // Nios_custom_instruction_master_translator:multi_ci_master_b -> Nios_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_c;             // Nios_custom_instruction_master_translator:multi_ci_master_c -> Nios_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_a;             // Nios_custom_instruction_master_translator:multi_ci_master_a -> Nios_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         nios_custom_instruction_master_translator_multi_ci_master_clk_en;        // Nios_custom_instruction_master_translator:multi_ci_master_clken -> Nios_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         nios_custom_instruction_master_translator_multi_ci_master_done;          // Nios_custom_instruction_master_multi_xconnect:ci_slave_done -> Nios_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios_custom_instruction_master_translator_multi_ci_master_n;             // Nios_custom_instruction_master_translator:multi_ci_master_n -> Nios_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         nios_custom_instruction_master_translator_multi_ci_master_writerc;       // Nios_custom_instruction_master_translator:multi_ci_master_writerc -> Nios_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios_custom_instruction_master_translator_multi_ci_master_clk;           // Nios_custom_instruction_master_translator:multi_ci_master_clk -> Nios_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios_custom_instruction_master_translator_multi_ci_master_reset_req;     // Nios_custom_instruction_master_translator:multi_ci_master_reset_req -> Nios_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios_custom_instruction_master_translator_multi_ci_master_start;         // Nios_custom_instruction_master_translator:multi_ci_master_start -> Nios_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_dataa;         // Nios_custom_instruction_master_translator:multi_ci_master_dataa -> Nios_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios_custom_instruction_master_translator_multi_ci_master_readra;        // Nios_custom_instruction_master_translator:multi_ci_master_readra -> Nios_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         nios_custom_instruction_master_translator_multi_ci_master_reset;         // Nios_custom_instruction_master_translator:multi_ci_master_reset -> Nios_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_datab;         // Nios_custom_instruction_master_translator:multi_ci_master_datab -> Nios_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         nios_custom_instruction_master_translator_multi_ci_master_readrb;        // Nios_custom_instruction_master_translator:multi_ci_master_readrb -> Nios_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_result;         // Nios_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Nios_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_b;              // Nios_custom_instruction_master_multi_xconnect:ci_master0_b -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_c;              // Nios_custom_instruction_master_multi_xconnect:ci_master0_c -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_done;           // Nios_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Nios_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // Nios_custom_instruction_master_multi_xconnect:ci_master0_clken -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_a;              // Nios_custom_instruction_master_multi_xconnect:ci_master0_a -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] nios_custom_instruction_master_multi_xconnect_ci_master0_n;              // Nios_custom_instruction_master_multi_xconnect:ci_master0_n -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // Nios_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // Nios_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_clk;            // Nios_custom_instruction_master_multi_xconnect:ci_master0_clk -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // Nios_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_start;          // Nios_custom_instruction_master_multi_xconnect:ci_master0_start -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // Nios_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_readra;         // Nios_custom_instruction_master_multi_xconnect:ci_master0_readra -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_reset;          // Nios_custom_instruction_master_multi_xconnect:ci_master0_reset -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_datab;          // Nios_custom_instruction_master_multi_xconnect:ci_master0_datab -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // Nios_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // Nios_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Nios_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_result; // LCD_0:result -> Nios_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_start;  // Nios_custom_instruction_master_multi_slave_translator0:ci_master_start -> LCD_0:start
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // Nios_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> LCD_0:dataa
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_done;   // LCD_0:done -> Nios_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // Nios_custom_instruction_master_multi_slave_translator0:ci_master_clken -> LCD_0:clk_en
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // Nios_custom_instruction_master_multi_slave_translator0:ci_master_reset -> LCD_0:reset
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // Nios_custom_instruction_master_multi_slave_translator0:ci_master_datab -> LCD_0:datab
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // Nios_custom_instruction_master_multi_slave_translator0:ci_master_clk -> LCD_0:clk
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                    // Jtag:av_waitrequest -> mm_interconnect_0:Jtag_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                      // mm_interconnect_0:Jtag_avalon_jtag_slave_writedata -> Jtag:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                        // mm_interconnect_0:Jtag_avalon_jtag_slave_address -> Jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                     // mm_interconnect_0:Jtag_avalon_jtag_slave_chipselect -> Jtag:av_chipselect
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                          // mm_interconnect_0:Jtag_avalon_jtag_slave_write -> Jtag:av_write_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                           // mm_interconnect_0:Jtag_avalon_jtag_slave_read -> Jtag:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                       // Jtag:av_readdata -> mm_interconnect_0:Jtag_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_led_3_s1_writedata;                                    // mm_interconnect_0:led_3_s1_writedata -> led_3:writedata
	wire   [1:0] mm_interconnect_0_led_3_s1_address;                                      // mm_interconnect_0:led_3_s1_address -> led_3:address
	wire         mm_interconnect_0_led_3_s1_chipselect;                                   // mm_interconnect_0:led_3_s1_chipselect -> led_3:chipselect
	wire         mm_interconnect_0_led_3_s1_write;                                        // mm_interconnect_0:led_3_s1_write -> led_3:write_n
	wire  [31:0] mm_interconnect_0_led_3_s1_readdata;                                     // led_3:readdata -> mm_interconnect_0:led_3_s1_readdata
	wire         nios_instruction_master_waitrequest;                                     // mm_interconnect_0:Nios_instruction_master_waitrequest -> Nios:i_waitrequest
	wire  [15:0] nios_instruction_master_address;                                         // Nios:i_address -> mm_interconnect_0:Nios_instruction_master_address
	wire         nios_instruction_master_read;                                            // Nios:i_read -> mm_interconnect_0:Nios_instruction_master_read
	wire  [31:0] nios_instruction_master_readdata;                                        // mm_interconnect_0:Nios_instruction_master_readdata -> Nios:i_readdata
	wire  [31:0] mm_interconnect_0_pushbutton_2_s1_writedata;                             // mm_interconnect_0:pushbutton_2_s1_writedata -> pushbutton_2:writedata
	wire   [1:0] mm_interconnect_0_pushbutton_2_s1_address;                               // mm_interconnect_0:pushbutton_2_s1_address -> pushbutton_2:address
	wire         mm_interconnect_0_pushbutton_2_s1_chipselect;                            // mm_interconnect_0:pushbutton_2_s1_chipselect -> pushbutton_2:chipselect
	wire         mm_interconnect_0_pushbutton_2_s1_write;                                 // mm_interconnect_0:pushbutton_2_s1_write -> pushbutton_2:write_n
	wire  [31:0] mm_interconnect_0_pushbutton_2_s1_readdata;                              // pushbutton_2:readdata -> mm_interconnect_0:pushbutton_2_s1_readdata
	wire   [1:0] mm_interconnect_0_dip_3_s1_address;                                      // mm_interconnect_0:dip_3_s1_address -> dip_3:address
	wire  [31:0] mm_interconnect_0_dip_3_s1_readdata;                                     // dip_3:readdata -> mm_interconnect_0:dip_3_s1_readdata
	wire  [31:0] mm_interconnect_0_led_1_s1_writedata;                                    // mm_interconnect_0:led_1_s1_writedata -> led_1:writedata
	wire   [1:0] mm_interconnect_0_led_1_s1_address;                                      // mm_interconnect_0:led_1_s1_address -> led_1:address
	wire         mm_interconnect_0_led_1_s1_chipselect;                                   // mm_interconnect_0:led_1_s1_chipselect -> led_1:chipselect
	wire         mm_interconnect_0_led_1_s1_write;                                        // mm_interconnect_0:led_1_s1_write -> led_1:write_n
	wire  [31:0] mm_interconnect_0_led_1_s1_readdata;                                     // led_1:readdata -> mm_interconnect_0:led_1_s1_readdata
	wire  [31:0] mm_interconnect_0_pushbutton_1_s1_writedata;                             // mm_interconnect_0:pushbutton_1_s1_writedata -> pushbutton_1:writedata
	wire   [1:0] mm_interconnect_0_pushbutton_1_s1_address;                               // mm_interconnect_0:pushbutton_1_s1_address -> pushbutton_1:address
	wire         mm_interconnect_0_pushbutton_1_s1_chipselect;                            // mm_interconnect_0:pushbutton_1_s1_chipselect -> pushbutton_1:chipselect
	wire         mm_interconnect_0_pushbutton_1_s1_write;                                 // mm_interconnect_0:pushbutton_1_s1_write -> pushbutton_1:write_n
	wire  [31:0] mm_interconnect_0_pushbutton_1_s1_readdata;                              // pushbutton_1:readdata -> mm_interconnect_0:pushbutton_1_s1_readdata
	wire   [1:0] mm_interconnect_0_dip_1_s1_address;                                      // mm_interconnect_0:dip_1_s1_address -> dip_1:address
	wire  [31:0] mm_interconnect_0_dip_1_s1_readdata;                                     // dip_1:readdata -> mm_interconnect_0:dip_1_s1_readdata
	wire  [31:0] mm_interconnect_0_led_2_s1_writedata;                                    // mm_interconnect_0:led_2_s1_writedata -> led_2:writedata
	wire   [1:0] mm_interconnect_0_led_2_s1_address;                                      // mm_interconnect_0:led_2_s1_address -> led_2:address
	wire         mm_interconnect_0_led_2_s1_chipselect;                                   // mm_interconnect_0:led_2_s1_chipselect -> led_2:chipselect
	wire         mm_interconnect_0_led_2_s1_write;                                        // mm_interconnect_0:led_2_s1_write -> led_2:write_n
	wire  [31:0] mm_interconnect_0_led_2_s1_readdata;                                     // led_2:readdata -> mm_interconnect_0:led_2_s1_readdata
	wire   [1:0] mm_interconnect_0_dip_0_s1_address;                                      // mm_interconnect_0:dip_0_s1_address -> dip_0:address
	wire  [31:0] mm_interconnect_0_dip_0_s1_readdata;                                     // dip_0:readdata -> mm_interconnect_0:dip_0_s1_readdata
	wire         mm_interconnect_0_nios_jtag_debug_module_waitrequest;                    // Nios:jtag_debug_module_waitrequest -> mm_interconnect_0:Nios_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios_jtag_debug_module_writedata;                      // mm_interconnect_0:Nios_jtag_debug_module_writedata -> Nios:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios_jtag_debug_module_address;                        // mm_interconnect_0:Nios_jtag_debug_module_address -> Nios:jtag_debug_module_address
	wire         mm_interconnect_0_nios_jtag_debug_module_write;                          // mm_interconnect_0:Nios_jtag_debug_module_write -> Nios:jtag_debug_module_write
	wire         mm_interconnect_0_nios_jtag_debug_module_read;                           // mm_interconnect_0:Nios_jtag_debug_module_read -> Nios:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios_jtag_debug_module_readdata;                       // Nios:jtag_debug_module_readdata -> mm_interconnect_0:Nios_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios_jtag_debug_module_debugaccess;                    // mm_interconnect_0:Nios_jtag_debug_module_debugaccess -> Nios:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios_jtag_debug_module_byteenable;                     // mm_interconnect_0:Nios_jtag_debug_module_byteenable -> Nios:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_led_5_s1_writedata;                                    // mm_interconnect_0:led_5_s1_writedata -> led_5:writedata
	wire   [1:0] mm_interconnect_0_led_5_s1_address;                                      // mm_interconnect_0:led_5_s1_address -> led_5:address
	wire         mm_interconnect_0_led_5_s1_chipselect;                                   // mm_interconnect_0:led_5_s1_chipselect -> led_5:chipselect
	wire         mm_interconnect_0_led_5_s1_write;                                        // mm_interconnect_0:led_5_s1_write -> led_5:write_n
	wire  [31:0] mm_interconnect_0_led_5_s1_readdata;                                     // led_5:readdata -> mm_interconnect_0:led_5_s1_readdata
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                                   // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire  [11:0] mm_interconnect_0_memory_s1_address;                                     // mm_interconnect_0:memory_s1_address -> memory:address
	wire         mm_interconnect_0_memory_s1_chipselect;                                  // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire         mm_interconnect_0_memory_s1_clken;                                       // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire         mm_interconnect_0_memory_s1_write;                                       // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                                    // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                                  // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         nios_data_master_waitrequest;                                            // mm_interconnect_0:Nios_data_master_waitrequest -> Nios:d_waitrequest
	wire  [31:0] nios_data_master_writedata;                                              // Nios:d_writedata -> mm_interconnect_0:Nios_data_master_writedata
	wire  [15:0] nios_data_master_address;                                                // Nios:d_address -> mm_interconnect_0:Nios_data_master_address
	wire         nios_data_master_write;                                                  // Nios:d_write -> mm_interconnect_0:Nios_data_master_write
	wire         nios_data_master_read;                                                   // Nios:d_read -> mm_interconnect_0:Nios_data_master_read
	wire  [31:0] nios_data_master_readdata;                                               // mm_interconnect_0:Nios_data_master_readdata -> Nios:d_readdata
	wire         nios_data_master_debugaccess;                                            // Nios:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:Nios_data_master_debugaccess
	wire   [3:0] nios_data_master_byteenable;                                             // Nios:d_byteenable -> mm_interconnect_0:Nios_data_master_byteenable
	wire   [1:0] mm_interconnect_0_dip_2_s1_address;                                      // mm_interconnect_0:dip_2_s1_address -> dip_2:address
	wire  [31:0] mm_interconnect_0_dip_2_s1_readdata;                                     // dip_2:readdata -> mm_interconnect_0:dip_2_s1_readdata
	wire  [31:0] mm_interconnect_0_led_4_s1_writedata;                                    // mm_interconnect_0:led_4_s1_writedata -> led_4:writedata
	wire   [1:0] mm_interconnect_0_led_4_s1_address;                                      // mm_interconnect_0:led_4_s1_address -> led_4:address
	wire         mm_interconnect_0_led_4_s1_chipselect;                                   // mm_interconnect_0:led_4_s1_chipselect -> led_4:chipselect
	wire         mm_interconnect_0_led_4_s1_write;                                        // mm_interconnect_0:led_4_s1_write -> led_4:write_n
	wire  [31:0] mm_interconnect_0_led_4_s1_readdata;                                     // led_4:readdata -> mm_interconnect_0:led_4_s1_readdata
	wire         mm_interconnect_0_eth_tse_0_control_port_waitrequest;                    // eth_tse_0:waitrequest -> mm_interconnect_0:eth_tse_0_control_port_waitrequest
	wire  [31:0] mm_interconnect_0_eth_tse_0_control_port_writedata;                      // mm_interconnect_0:eth_tse_0_control_port_writedata -> eth_tse_0:writedata
	wire   [7:0] mm_interconnect_0_eth_tse_0_control_port_address;                        // mm_interconnect_0:eth_tse_0_control_port_address -> eth_tse_0:address
	wire         mm_interconnect_0_eth_tse_0_control_port_write;                          // mm_interconnect_0:eth_tse_0_control_port_write -> eth_tse_0:write
	wire         mm_interconnect_0_eth_tse_0_control_port_read;                           // mm_interconnect_0:eth_tse_0_control_port_read -> eth_tse_0:read
	wire  [31:0] mm_interconnect_0_eth_tse_0_control_port_readdata;                       // eth_tse_0:readdata -> mm_interconnect_0:eth_tse_0_control_port_readdata
	wire         irq_mapper_receiver0_irq;                                                // Jtag:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_d_irq_irq;                                                          // irq_mapper:sender_irq -> Nios:d_irq
	wire         eth_tse_0_receive_endofpacket;                                           // eth_tse_0:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire         eth_tse_0_receive_valid;                                                 // eth_tse_0:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire         eth_tse_0_receive_startofpacket;                                         // eth_tse_0:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire   [5:0] eth_tse_0_receive_error;                                                 // eth_tse_0:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] eth_tse_0_receive_empty;                                                 // eth_tse_0:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire  [31:0] eth_tse_0_receive_data;                                                  // eth_tse_0:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         eth_tse_0_receive_ready;                                                 // avalon_st_adapter:in_0_ready -> eth_tse_0:ff_rx_rdy
	wire         avalon_st_adapter_out_0_endofpacket;                                     // avalon_st_adapter:out_0_endofpacket -> eth_tse_0:ff_tx_eop
	wire         avalon_st_adapter_out_0_valid;                                           // avalon_st_adapter:out_0_valid -> eth_tse_0:ff_tx_wren
	wire         avalon_st_adapter_out_0_startofpacket;                                   // avalon_st_adapter:out_0_startofpacket -> eth_tse_0:ff_tx_sop
	wire         avalon_st_adapter_out_0_error;                                           // avalon_st_adapter:out_0_error -> eth_tse_0:ff_tx_err
	wire   [1:0] avalon_st_adapter_out_0_empty;                                           // avalon_st_adapter:out_0_empty -> eth_tse_0:ff_tx_mod
	wire  [31:0] avalon_st_adapter_out_0_data;                                            // avalon_st_adapter:out_0_data -> eth_tse_0:ff_tx_data
	wire         avalon_st_adapter_out_0_ready;                                           // eth_tse_0:ff_tx_rdy -> avalon_st_adapter:out_0_ready
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [Jtag:rst_n, Nios:reset_n, dip_0:reset_n, dip_1:reset_n, dip_2:reset_n, dip_3:reset_n, irq_mapper:reset, led_1:reset_n, led_2:reset_n, led_3:reset_n, led_4:reset_n, led_5:reset_n, memory:reset, mm_interconnect_0:Nios_reset_n_reset_bridge_in_reset_reset, pushbutton_1:reset_n, pushbutton_2:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [Nios:reset_req, memory:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, eth_tse_0:reset, mm_interconnect_0:eth_tse_0_reset_connection_reset_bridge_in_reset_reset]

	Nios_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)      //       .reset_req
	);

	Nios_Nios nios (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (nios_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios_data_master_read),                                //                          .read
		.d_readdata                            (nios_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios_data_master_write),                               //                          .write
		.d_writedata                           (nios_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios_instruction_master_read),                         //                          .read
		.i_readdata                            (nios_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_multi_done                       (nios_custom_instruction_master_done),                  // custom_instruction_master.done
		.E_ci_multi_clk_en                     (nios_custom_instruction_master_clk_en),                //                          .clk_en
		.E_ci_multi_start                      (nios_custom_instruction_master_start),                 //                          .start
		.E_ci_result                           (nios_custom_instruction_master_result),                //                          .result
		.D_ci_a                                (nios_custom_instruction_master_a),                     //                          .a
		.D_ci_b                                (nios_custom_instruction_master_b),                     //                          .b
		.D_ci_c                                (nios_custom_instruction_master_c),                     //                          .c
		.D_ci_n                                (nios_custom_instruction_master_n),                     //                          .n
		.D_ci_readra                           (nios_custom_instruction_master_readra),                //                          .readra
		.D_ci_readrb                           (nios_custom_instruction_master_readrb),                //                          .readrb
		.D_ci_writerc                          (nios_custom_instruction_master_writerc),               //                          .writerc
		.E_ci_dataa                            (nios_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_datab                            (nios_custom_instruction_master_datab),                 //                          .datab
		.E_ci_multi_clock                      (nios_custom_instruction_master_clk),                   //                          .clk
		.E_ci_multi_reset                      (nios_custom_instruction_master_reset),                 //                          .reset
		.E_ci_multi_reset_req                  (nios_custom_instruction_master_reset_req)              //                          .reset_req
	);

	Nios_Jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	Nios_pushbutton_2 pushbutton_2 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_pushbutton_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pushbutton_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pushbutton_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pushbutton_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pushbutton_2_s1_readdata),   //                    .readdata
		.in_port    (pushbutton2_external_connection_export)        // external_connection.export
	);

	Nios_led_1 led_1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_1_s1_readdata),   //                    .readdata
		.out_port   (led_1_external_connection_export)       // external_connection.export
	);

	Nios_led_1 led_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_2_s1_readdata),   //                    .readdata
		.out_port   (led_2_external_connection_export)       // external_connection.export
	);

	Nios_led_1 led_3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_3_s1_readdata),   //                    .readdata
		.out_port   (led_3_external_connection_export)       // external_connection.export
	);

	Nios_led_1 led_4 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_4_s1_readdata),   //                    .readdata
		.out_port   (led_4_external_connection_export)       // external_connection.export
	);

	Nios_led_1 led_5 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_5_s1_readdata),   //                    .readdata
		.out_port   (led_5_external_connection_export)       // external_connection.export
	);

	Nios_pushbutton_2 pushbutton_1 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_pushbutton_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pushbutton_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pushbutton_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pushbutton_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pushbutton_1_s1_readdata),   //                    .readdata
		.in_port    (pushbutton_1_external_connection_export)       // external_connection.export
	);

	Nios_dip_0 dip_0 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_dip_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dip_0_s1_readdata), //                    .readdata
		.in_port  (dip_0_external_connection_export)     // external_connection.export
	);

	Nios_dip_0 dip_1 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_dip_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dip_1_s1_readdata), //                    .readdata
		.in_port  (dip_1_external_connection_export)     // external_connection.export
	);

	Nios_dip_0 dip_2 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_dip_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dip_2_s1_readdata), //                    .readdata
		.in_port  (dip_2_external_connection_export)     // external_connection.export
	);

	Nios_dip_0 dip_3 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_dip_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dip_3_s1_readdata), //                    .readdata
		.in_port  (dip_3_external_connection_export)     // external_connection.export
	);

	lcd_driver lcd_0 (
		.rs     (lcd_0_conduit_end_rs),                                                    //                     conduit_end.export
		.rw     (lcd_0_conduit_end_rw),                                                    //                                .export
		.en     (lcd_0_conduit_end_en),                                                    //                                .export
		.db     (lcd_0_conduit_end_db),                                                    //                                .export
		.dataa  (nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave_3.dataa
		.datab  (nios_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                                .datab
		.result (nios_custom_instruction_master_multi_slave_translator0_ci_master_result), //                                .result
		.clk    (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                                .clk
		.clk_en (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                                .clk_en
		.start  (nios_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                                .start
		.reset  (nios_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                                .reset
		.done   (nios_custom_instruction_master_multi_slave_translator0_ci_master_done)    //                                .done
	);

	Nios_eth_tse_0 eth_tse_0 (
		.clk           (clk_clk),                                              // control_port_clock_connection.clk
		.reset         (rst_controller_001_reset_out_reset),                   //              reset_connection.reset
		.address       (mm_interconnect_0_eth_tse_0_control_port_address),     //                  control_port.address
		.readdata      (mm_interconnect_0_eth_tse_0_control_port_readdata),    //                              .readdata
		.read          (mm_interconnect_0_eth_tse_0_control_port_read),        //                              .read
		.writedata     (mm_interconnect_0_eth_tse_0_control_port_writedata),   //                              .writedata
		.write         (mm_interconnect_0_eth_tse_0_control_port_write),       //                              .write
		.waitrequest   (mm_interconnect_0_eth_tse_0_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (clk_clk),                                              //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (clk_clk),                                              //   pcs_mac_rx_clock_connection.clk
		.set_10        (eth_tse_0_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (eth_tse_0_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (eth_tse_0_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (eth_tse_0_mac_status_connection_ena_10),               //                              .ena_10
		.gm_rx_d       (eth_tse_0_mac_gmii_connection_gmii_rx_d),              //           mac_gmii_connection.gmii_rx_d
		.gm_rx_dv      (eth_tse_0_mac_gmii_connection_gmii_rx_dv),             //                              .gmii_rx_dv
		.gm_rx_err     (eth_tse_0_mac_gmii_connection_gmii_rx_err),            //                              .gmii_rx_err
		.gm_tx_d       (eth_tse_0_mac_gmii_connection_gmii_tx_d),              //                              .gmii_tx_d
		.gm_tx_en      (eth_tse_0_mac_gmii_connection_gmii_tx_en),             //                              .gmii_tx_en
		.gm_tx_err     (eth_tse_0_mac_gmii_connection_gmii_tx_err),            //                              .gmii_tx_err
		.m_rx_d        (eth_tse_0_mac_mii_connection_mii_rx_d),                //            mac_mii_connection.mii_rx_d
		.m_rx_en       (eth_tse_0_mac_mii_connection_mii_rx_dv),               //                              .mii_rx_dv
		.m_rx_err      (eth_tse_0_mac_mii_connection_mii_rx_err),              //                              .mii_rx_err
		.m_tx_d        (eth_tse_0_mac_mii_connection_mii_tx_d),                //                              .mii_tx_d
		.m_tx_en       (eth_tse_0_mac_mii_connection_mii_tx_en),               //                              .mii_tx_en
		.m_tx_err      (eth_tse_0_mac_mii_connection_mii_tx_err),              //                              .mii_tx_err
		.m_rx_crs      (eth_tse_0_mac_mii_connection_mii_crs),                 //                              .mii_crs
		.m_rx_col      (eth_tse_0_mac_mii_connection_mii_col),                 //                              .mii_col
		.ff_rx_clk     (clk_clk),                                              //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                              //     transmit_clock_connection.clk
		.ff_rx_data    (eth_tse_0_receive_data),                               //                       receive.data
		.ff_rx_eop     (eth_tse_0_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (eth_tse_0_receive_error),                              //                              .error
		.ff_rx_mod     (eth_tse_0_receive_empty),                              //                              .empty
		.ff_rx_rdy     (eth_tse_0_receive_ready),                              //                              .ready
		.ff_rx_sop     (eth_tse_0_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (eth_tse_0_receive_valid),                              //                              .valid
		.ff_tx_data    (avalon_st_adapter_out_0_data),                         //                      transmit.data
		.ff_tx_eop     (avalon_st_adapter_out_0_endofpacket),                  //                              .endofpacket
		.ff_tx_err     (avalon_st_adapter_out_0_error),                        //                              .error
		.ff_tx_mod     (avalon_st_adapter_out_0_empty),                        //                              .empty
		.ff_tx_rdy     (avalon_st_adapter_out_0_ready),                        //                              .ready
		.ff_tx_sop     (avalon_st_adapter_out_0_startofpacket),                //                              .startofpacket
		.ff_tx_wren    (avalon_st_adapter_out_0_valid),                        //                              .valid
		.magic_wakeup  (eth_tse_0_mac_misc_connection_magic_wakeup),           //           mac_misc_connection.magic_wakeup
		.magic_sleep_n (eth_tse_0_mac_misc_connection_magic_sleep_n),          //                              .magic_sleep_n
		.ff_tx_crc_fwd (eth_tse_0_mac_misc_connection_ff_tx_crc_fwd),          //                              .ff_tx_crc_fwd
		.ff_tx_septy   (eth_tse_0_mac_misc_connection_ff_tx_septy),            //                              .ff_tx_septy
		.tx_ff_uflow   (eth_tse_0_mac_misc_connection_tx_ff_uflow),            //                              .tx_ff_uflow
		.ff_tx_a_full  (eth_tse_0_mac_misc_connection_ff_tx_a_full),           //                              .ff_tx_a_full
		.ff_tx_a_empty (eth_tse_0_mac_misc_connection_ff_tx_a_empty),          //                              .ff_tx_a_empty
		.rx_err_stat   (eth_tse_0_mac_misc_connection_rx_err_stat),            //                              .rx_err_stat
		.rx_frm_type   (eth_tse_0_mac_misc_connection_rx_frm_type),            //                              .rx_frm_type
		.ff_rx_dsav    (eth_tse_0_mac_misc_connection_ff_rx_dsav),             //                              .ff_rx_dsav
		.ff_rx_a_full  (eth_tse_0_mac_misc_connection_ff_rx_a_full),           //                              .ff_rx_a_full
		.ff_rx_a_empty (eth_tse_0_mac_misc_connection_ff_rx_a_empty)           //                              .ff_rx_a_empty
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios_custom_instruction_master_translator (
		.ci_slave_dataa            (nios_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (),                                                                    //                .ipending
		.ci_slave_estatus          (),                                                                    //                .estatus
		.ci_slave_multi_clk        (nios_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                    //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                    //                .datab
		.comb_ci_master_result     (),                                                                    //                .result
		.comb_ci_master_n          (),                                                                    //                .n
		.comb_ci_master_readra     (),                                                                    //                .readra
		.comb_ci_master_readrb     (),                                                                    //                .readrb
		.comb_ci_master_writerc    (),                                                                    //                .writerc
		.comb_ci_master_a          (),                                                                    //                .a
		.comb_ci_master_b          (),                                                                    //                .b
		.comb_ci_master_c          (),                                                                    //                .c
		.comb_ci_master_ipending   (),                                                                    //                .ipending
		.comb_ci_master_estatus    (),                                                                    //                .estatus
		.multi_ci_master_clk       (nios_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                //     (terminated)
		.ci_slave_multi_result     (),                                                                    //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                         //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                            //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                            //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                             //     (terminated)
	);

	Nios_Nios_custom_instruction_master_multi_xconnect nios_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                    //           .ipending
		.ci_slave_estatus     (),                                                                    //           .estatus
		.ci_slave_clk         (nios_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_clk       (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_n         (),                                                                        // (terminated)
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_reset_req ()                                                                         // (terminated)
	);

	Nios_mm_interconnect_0 mm_interconnect_0 (
		.Clk_clk_clk                                            (clk_clk),                                              //                                          Clk_clk.clk
		.eth_tse_0_reset_connection_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                   // eth_tse_0_reset_connection_reset_bridge_in_reset.reset
		.Nios_reset_n_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                       //               Nios_reset_n_reset_bridge_in_reset.reset
		.Nios_data_master_address                               (nios_data_master_address),                             //                                 Nios_data_master.address
		.Nios_data_master_waitrequest                           (nios_data_master_waitrequest),                         //                                                 .waitrequest
		.Nios_data_master_byteenable                            (nios_data_master_byteenable),                          //                                                 .byteenable
		.Nios_data_master_read                                  (nios_data_master_read),                                //                                                 .read
		.Nios_data_master_readdata                              (nios_data_master_readdata),                            //                                                 .readdata
		.Nios_data_master_write                                 (nios_data_master_write),                               //                                                 .write
		.Nios_data_master_writedata                             (nios_data_master_writedata),                           //                                                 .writedata
		.Nios_data_master_debugaccess                           (nios_data_master_debugaccess),                         //                                                 .debugaccess
		.Nios_instruction_master_address                        (nios_instruction_master_address),                      //                          Nios_instruction_master.address
		.Nios_instruction_master_waitrequest                    (nios_instruction_master_waitrequest),                  //                                                 .waitrequest
		.Nios_instruction_master_read                           (nios_instruction_master_read),                         //                                                 .read
		.Nios_instruction_master_readdata                       (nios_instruction_master_readdata),                     //                                                 .readdata
		.dip_0_s1_address                                       (mm_interconnect_0_dip_0_s1_address),                   //                                         dip_0_s1.address
		.dip_0_s1_readdata                                      (mm_interconnect_0_dip_0_s1_readdata),                  //                                                 .readdata
		.dip_1_s1_address                                       (mm_interconnect_0_dip_1_s1_address),                   //                                         dip_1_s1.address
		.dip_1_s1_readdata                                      (mm_interconnect_0_dip_1_s1_readdata),                  //                                                 .readdata
		.dip_2_s1_address                                       (mm_interconnect_0_dip_2_s1_address),                   //                                         dip_2_s1.address
		.dip_2_s1_readdata                                      (mm_interconnect_0_dip_2_s1_readdata),                  //                                                 .readdata
		.dip_3_s1_address                                       (mm_interconnect_0_dip_3_s1_address),                   //                                         dip_3_s1.address
		.dip_3_s1_readdata                                      (mm_interconnect_0_dip_3_s1_readdata),                  //                                                 .readdata
		.eth_tse_0_control_port_address                         (mm_interconnect_0_eth_tse_0_control_port_address),     //                           eth_tse_0_control_port.address
		.eth_tse_0_control_port_write                           (mm_interconnect_0_eth_tse_0_control_port_write),       //                                                 .write
		.eth_tse_0_control_port_read                            (mm_interconnect_0_eth_tse_0_control_port_read),        //                                                 .read
		.eth_tse_0_control_port_readdata                        (mm_interconnect_0_eth_tse_0_control_port_readdata),    //                                                 .readdata
		.eth_tse_0_control_port_writedata                       (mm_interconnect_0_eth_tse_0_control_port_writedata),   //                                                 .writedata
		.eth_tse_0_control_port_waitrequest                     (mm_interconnect_0_eth_tse_0_control_port_waitrequest), //                                                 .waitrequest
		.Jtag_avalon_jtag_slave_address                         (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                           Jtag_avalon_jtag_slave.address
		.Jtag_avalon_jtag_slave_write                           (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                                 .write
		.Jtag_avalon_jtag_slave_read                            (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                                 .read
		.Jtag_avalon_jtag_slave_readdata                        (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                                 .readdata
		.Jtag_avalon_jtag_slave_writedata                       (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                                 .writedata
		.Jtag_avalon_jtag_slave_waitrequest                     (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                                 .waitrequest
		.Jtag_avalon_jtag_slave_chipselect                      (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                                 .chipselect
		.led_1_s1_address                                       (mm_interconnect_0_led_1_s1_address),                   //                                         led_1_s1.address
		.led_1_s1_write                                         (mm_interconnect_0_led_1_s1_write),                     //                                                 .write
		.led_1_s1_readdata                                      (mm_interconnect_0_led_1_s1_readdata),                  //                                                 .readdata
		.led_1_s1_writedata                                     (mm_interconnect_0_led_1_s1_writedata),                 //                                                 .writedata
		.led_1_s1_chipselect                                    (mm_interconnect_0_led_1_s1_chipselect),                //                                                 .chipselect
		.led_2_s1_address                                       (mm_interconnect_0_led_2_s1_address),                   //                                         led_2_s1.address
		.led_2_s1_write                                         (mm_interconnect_0_led_2_s1_write),                     //                                                 .write
		.led_2_s1_readdata                                      (mm_interconnect_0_led_2_s1_readdata),                  //                                                 .readdata
		.led_2_s1_writedata                                     (mm_interconnect_0_led_2_s1_writedata),                 //                                                 .writedata
		.led_2_s1_chipselect                                    (mm_interconnect_0_led_2_s1_chipselect),                //                                                 .chipselect
		.led_3_s1_address                                       (mm_interconnect_0_led_3_s1_address),                   //                                         led_3_s1.address
		.led_3_s1_write                                         (mm_interconnect_0_led_3_s1_write),                     //                                                 .write
		.led_3_s1_readdata                                      (mm_interconnect_0_led_3_s1_readdata),                  //                                                 .readdata
		.led_3_s1_writedata                                     (mm_interconnect_0_led_3_s1_writedata),                 //                                                 .writedata
		.led_3_s1_chipselect                                    (mm_interconnect_0_led_3_s1_chipselect),                //                                                 .chipselect
		.led_4_s1_address                                       (mm_interconnect_0_led_4_s1_address),                   //                                         led_4_s1.address
		.led_4_s1_write                                         (mm_interconnect_0_led_4_s1_write),                     //                                                 .write
		.led_4_s1_readdata                                      (mm_interconnect_0_led_4_s1_readdata),                  //                                                 .readdata
		.led_4_s1_writedata                                     (mm_interconnect_0_led_4_s1_writedata),                 //                                                 .writedata
		.led_4_s1_chipselect                                    (mm_interconnect_0_led_4_s1_chipselect),                //                                                 .chipselect
		.led_5_s1_address                                       (mm_interconnect_0_led_5_s1_address),                   //                                         led_5_s1.address
		.led_5_s1_write                                         (mm_interconnect_0_led_5_s1_write),                     //                                                 .write
		.led_5_s1_readdata                                      (mm_interconnect_0_led_5_s1_readdata),                  //                                                 .readdata
		.led_5_s1_writedata                                     (mm_interconnect_0_led_5_s1_writedata),                 //                                                 .writedata
		.led_5_s1_chipselect                                    (mm_interconnect_0_led_5_s1_chipselect),                //                                                 .chipselect
		.memory_s1_address                                      (mm_interconnect_0_memory_s1_address),                  //                                        memory_s1.address
		.memory_s1_write                                        (mm_interconnect_0_memory_s1_write),                    //                                                 .write
		.memory_s1_readdata                                     (mm_interconnect_0_memory_s1_readdata),                 //                                                 .readdata
		.memory_s1_writedata                                    (mm_interconnect_0_memory_s1_writedata),                //                                                 .writedata
		.memory_s1_byteenable                                   (mm_interconnect_0_memory_s1_byteenable),               //                                                 .byteenable
		.memory_s1_chipselect                                   (mm_interconnect_0_memory_s1_chipselect),               //                                                 .chipselect
		.memory_s1_clken                                        (mm_interconnect_0_memory_s1_clken),                    //                                                 .clken
		.Nios_jtag_debug_module_address                         (mm_interconnect_0_nios_jtag_debug_module_address),     //                           Nios_jtag_debug_module.address
		.Nios_jtag_debug_module_write                           (mm_interconnect_0_nios_jtag_debug_module_write),       //                                                 .write
		.Nios_jtag_debug_module_read                            (mm_interconnect_0_nios_jtag_debug_module_read),        //                                                 .read
		.Nios_jtag_debug_module_readdata                        (mm_interconnect_0_nios_jtag_debug_module_readdata),    //                                                 .readdata
		.Nios_jtag_debug_module_writedata                       (mm_interconnect_0_nios_jtag_debug_module_writedata),   //                                                 .writedata
		.Nios_jtag_debug_module_byteenable                      (mm_interconnect_0_nios_jtag_debug_module_byteenable),  //                                                 .byteenable
		.Nios_jtag_debug_module_waitrequest                     (mm_interconnect_0_nios_jtag_debug_module_waitrequest), //                                                 .waitrequest
		.Nios_jtag_debug_module_debugaccess                     (mm_interconnect_0_nios_jtag_debug_module_debugaccess), //                                                 .debugaccess
		.pushbutton_1_s1_address                                (mm_interconnect_0_pushbutton_1_s1_address),            //                                  pushbutton_1_s1.address
		.pushbutton_1_s1_write                                  (mm_interconnect_0_pushbutton_1_s1_write),              //                                                 .write
		.pushbutton_1_s1_readdata                               (mm_interconnect_0_pushbutton_1_s1_readdata),           //                                                 .readdata
		.pushbutton_1_s1_writedata                              (mm_interconnect_0_pushbutton_1_s1_writedata),          //                                                 .writedata
		.pushbutton_1_s1_chipselect                             (mm_interconnect_0_pushbutton_1_s1_chipselect),         //                                                 .chipselect
		.pushbutton_2_s1_address                                (mm_interconnect_0_pushbutton_2_s1_address),            //                                  pushbutton_2_s1.address
		.pushbutton_2_s1_write                                  (mm_interconnect_0_pushbutton_2_s1_write),              //                                                 .write
		.pushbutton_2_s1_readdata                               (mm_interconnect_0_pushbutton_2_s1_readdata),           //                                                 .readdata
		.pushbutton_2_s1_writedata                              (mm_interconnect_0_pushbutton_2_s1_writedata),          //                                                 .writedata
		.pushbutton_2_s1_chipselect                             (mm_interconnect_0_pushbutton_2_s1_chipselect)          //                                                 .chipselect
	);

	Nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_d_irq_irq)                  //    sender.irq
	);

	Nios_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),    // in_rst_0.reset
		.in_0_ready          (eth_tse_0_receive_ready),               //     in_0.ready
		.in_0_valid          (eth_tse_0_receive_valid),               //         .valid
		.in_0_data           (eth_tse_0_receive_data),                //         .data
		.in_0_startofpacket  (eth_tse_0_receive_startofpacket),       //         .startofpacket
		.in_0_endofpacket    (eth_tse_0_receive_endofpacket),         //         .endofpacket
		.in_0_empty          (eth_tse_0_receive_empty),               //         .empty
		.in_0_error          (eth_tse_0_receive_error),               //         .error
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //    out_0.ready
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_data          (avalon_st_adapter_out_0_data),          //         .data
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (nios_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios_jtag_debug_module_reset_reset), // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
